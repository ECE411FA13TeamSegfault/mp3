CONFIGURATION Memory_untitled_config OF Memory IS
   FOR untitled
   END FOR;
END Memory_untitled_config;