CONFIGURATION BRadd_untitled_config OF BRadd IS
   FOR untitled
   END FOR;
END BRadd_untitled_config;