--
-- VHDL Architecture ece411.SEXT4.untitled
--
-- Created:
--          by - chng2.ews (linux-a2.ews.illinois.edu)
--          at - 11:36:57 09/13/13
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY SEXT4 IS
   PORT( 
      clk : IN     std_logic
   );

-- Declarations

END SEXT4 ;

--
ARCHITECTURE untitled OF SEXT4 IS
BEGIN
END ARCHITECTURE untitled;

