CONFIGURATION AND2_UNTITLED_config OF AND2 IS
   FOR UNTITLED
   END FOR;
END AND2_UNTITLED_config;