CONFIGURATION NAND3_UNTITLED_config OF NAND3 IS
   FOR UNTITLED
   END FOR;
END NAND3_UNTITLED_config;