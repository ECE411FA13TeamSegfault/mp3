--
-- VHDL Architecture ece411.PredictArray.untitled
--
-- Created:
--          by - chao16.ews (gelib-057-38.ews.illinois.edu)
--          at - 00:52:15 09/19/13
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY PredictArray IS
   PORT( 
      Input     : IN     std_logic_vector(1 downto 0);
      WriteEN   : IN     std_logic;
      Index     : IN     LC3B_C_INDEX;
      RESET_L   : IN     std_logic;
      Output    : OUT    std_logic_vector(1 downto 0);
      clk       : IN     std_logic
   );

-- Declarations

END PredictArray ;

--
ARCHITECTURE untitled OF PredictArray IS
  TYPE PredictArray IS array (7 downto 0) of std_logic_vector(1 downto 0);
  SIGNAL Predict : PredictArray;
BEGIN
  ------------------------------------------------------------------
  ReadFromPredictArray: PROCESS (Predict, Index)
  ------------------------------------------------------------------
  VARIABLE PredictIndex : integer;
  BEGIN
    PredictIndex := to_integer(unsigned(Index));
    Output <= Predict(PredictIndex) after DELAY_256B;
  END PROCESS ReadFromPredictArray;
  ------------------------------------------------------------------
  WriteToPredictArray: PROCESS (clk, RESET_L, Index, WriteEN, Input)
  ------------------------------------------------------------------
  VARIABLE PredictIndex : integer;
  BEGIN
    PredictIndex := to_integer(unsigned(Index));
    IF RESET_L = '0' THEN
      Predict(0) <= (OTHERS => 'X');
      Predict(1) <= (OTHERS => 'X');
      Predict(2) <= (OTHERS => 'X');
      Predict(3) <= (OTHERS => 'X');
      Predict(4) <= (OTHERS => 'X');
      Predict(5) <= (OTHERS => 'X');
      Predict(6) <= (OTHERS => 'X');
      Predict(7) <= (OTHERS => 'X');
    END IF;
    if (clk'event and (clk = '1') and (clk'last_value = '0')) then
      IF (WriteEN = '1') THEN
        Predict(PredictIndex) <= Input;
      END IF;
    end if;
  END PROCESS WriteToPredictArray;
END ARCHITECTURE untitled;

