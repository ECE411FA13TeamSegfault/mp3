CONFIGURATION NOT1_UNTITLED_config OF NOT1 IS
   FOR UNTITLED
   END FOR;
END NOT1_UNTITLED_config;