CONFIGURATION OR2_UNTITLED_config OF OR2 IS
   FOR UNTITLED
   END FOR;
END OR2_UNTITLED_config;