CONFIGURATION CLKgen_untitled_config OF CLKgen IS
   FOR untitled
   END FOR;
END CLKgen_untitled_config;