CONFIGURATION MUX2_1_UNTITLED_config OF MUX2_1 IS
   FOR UNTITLED
   END FOR;
END MUX2_1_UNTITLED_config;