CONFIGURATION NAND2_UNTITLED_config OF NAND2 IS
   FOR UNTITLED
   END FOR;
END NAND2_UNTITLED_config;