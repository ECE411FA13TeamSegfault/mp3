--
-- VHDL Architecture ece411.DEMUX2_16.untitled
--
-- Created:
--          by - chao16.ews (dcl-l520-09.ews.illinois.edu)
--          at - 18:28:57 11/14/13
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY DEMUX2_128 IS
   PORT( 
      F   : IN     LC3B_OWORD;
      Sel : IN     std_logic;
      A   : OUT    LC3B_OWORD;
      B   : OUT    LC3B_OWORD
   );

-- Declarations

END DEMUX2_128 ;

--
ARCHITECTURE untitled OF DEMUX2_128 IS
BEGIN
	DEMUX2_128: PROCESS(F, SEL)
	BEGIN
		CASE SEL IS
		WHEN '0' =>
			A <= F AFTER DELAY_MUX2;
			B <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" AFTER DELAY_MUX2;
		WHEN '1' =>
			B <= F AFTER DELAY_MUX2;
			A <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" AFTER DELAY_MUX2;
		WHEN OTHERS =>
			A <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" AFTER DELAY_MUX2;
			B <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" AFTER DELAY_MUX2;
		END CASE;
	END PROCESS DEMUX2_128;
END ARCHITECTURE untitled;

